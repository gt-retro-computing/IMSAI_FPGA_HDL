module uart_device_tb;

    reg reset = 1;
    
endmodule