
module uart_debug (
	source,
	probe);	

	output	[9:0]	source;
	input	[0:0]	probe;
endmodule
